
module Not(
	// Input signals
	input wire a,	
	// Output signals
	output wire b	
);
	assign b = ~a;

endmodule





